library verilog;
use verilog.vl_types.all;
entity somador8bits_vlg_vec_tst is
end somador8bits_vlg_vec_tst;
