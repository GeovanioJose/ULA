library verilog;
use verilog.vl_types.all;
entity AxorB8bits_vlg_vec_tst is
end AxorB8bits_vlg_vec_tst;
