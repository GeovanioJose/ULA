library verilog;
use verilog.vl_types.all;
entity AxnorB8bits_vlg_vec_tst is
end AxnorB8bits_vlg_vec_tst;
