library verilog;
use verilog.vl_types.all;
entity AxnorB8bits_vlg_check_tst is
    port(
        S               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end AxnorB8bits_vlg_check_tst;
